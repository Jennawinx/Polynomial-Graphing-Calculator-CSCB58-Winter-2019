module Hex_Display(IN, OUT);
    input [4:0] IN;
	output reg [6:0] OUT;

	always @(*)
	begin
		case(IN[4:0])
			5'b00000: OUT = 7'b1000000;	// 0
			5'b00001: OUT = 7'b1111001;	// 1
			5'b00010: OUT = 7'b0100100;	// 2
			5'b00011: OUT = 7'b0110000; // 3
			5'b00100: OUT = 7'b0011001; // 4
			5'b00101: OUT = 7'b0010010; // 5
			5'b00110: OUT = 7'b0000010; // 6
			5'b00111: OUT = 7'b1111000; // 7
			5'b01000: OUT = 7'b0000000; // 8
			5'b01001: OUT = 7'b0011000; // 9
			5'b01010: OUT = 7'b0001000; // A
			5'b01011: OUT = 7'b0000011; // b
			5'b01100: OUT = 7'b1000110; // C
			5'b01101: OUT = 7'b0100001; // d
			5'b01110: OUT = 7'b0000110; // E
			5'b01111: OUT = 7'b0001110; // F
			5'b10000: OUT = 7'b0101011;	// n
			5'b10001: OUT = 7'b0111111;	// -
			5'b10010: OUT = 7'b1000111;	// L
			5'b10011: OUT = 7'b0001100;	// p
			5'b10100: OUT = 7'b0010000; // g
			5'b10101: OUT = 7'b1001000;	// N
			default: OUT = 7'b1111111; // Blank
		endcase

	end

endmodule